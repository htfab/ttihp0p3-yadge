VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_htfab_yadge
  CLASS BLOCK ;
  FOREIGN tt_um_htfab_yadge ;
  ORIGIN 0.000 0.000 ;
  SIZE 202.080 BY 154.980 ;
  PIN clk
    PORT
      LAYER Metal5 ;
        RECT 187.050 153.980 187.350 154.980 ;
    END
  END clk
  PIN ena
    PORT
      LAYER Metal5 ;
        RECT 190.890 153.980 191.190 154.980 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER Metal5 ;
        RECT 183.210 153.980 183.510 154.980 ;
    END
  END rst_n
  PIN ui_in[0]
    PORT
      LAYER Metal5 ;
        RECT 179.370 153.980 179.670 154.980 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER Metal5 ;
        RECT 175.530 153.980 175.830 154.980 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER Metal5 ;
        RECT 171.690 153.980 171.990 154.980 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER Metal5 ;
        RECT 167.850 153.980 168.150 154.980 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER Metal5 ;
        RECT 164.010 153.980 164.310 154.980 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER Metal5 ;
        RECT 160.170 153.980 160.470 154.980 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER Metal5 ;
        RECT 156.330 153.980 156.630 154.980 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER Metal5 ;
        RECT 152.490 153.980 152.790 154.980 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER Metal5 ;
        RECT 148.650 153.980 148.950 154.980 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER Metal5 ;
        RECT 144.810 153.980 145.110 154.980 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER Metal5 ;
        RECT 140.970 153.980 141.270 154.980 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER Metal5 ;
        RECT 137.130 153.980 137.430 154.980 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER Metal5 ;
        RECT 133.290 153.980 133.590 154.980 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER Metal5 ;
        RECT 129.450 153.980 129.750 154.980 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER Metal5 ;
        RECT 125.610 153.980 125.910 154.980 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER Metal5 ;
        RECT 121.770 153.980 122.070 154.980 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER Metal5 ;
        RECT 56.490 153.980 56.790 154.980 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER Metal5 ;
        RECT 52.650 153.980 52.950 154.980 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    PORT
      LAYER Metal5 ;
        RECT 48.810 153.980 49.110 154.980 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER Metal5 ;
        RECT 44.970 153.980 45.270 154.980 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER Metal5 ;
        RECT 41.130 153.980 41.430 154.980 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER Metal5 ;
        RECT 37.290 153.980 37.590 154.980 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER Metal5 ;
        RECT 33.450 153.980 33.750 154.980 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER Metal5 ;
        RECT 29.610 153.980 29.910 154.980 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER Metal5 ;
        RECT 87.210 153.980 87.510 154.980 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER Metal5 ;
        RECT 83.370 153.980 83.670 154.980 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER Metal5 ;
        RECT 79.530 153.980 79.830 154.980 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER Metal5 ;
        RECT 75.690 153.980 75.990 154.980 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    PORT
      LAYER Metal5 ;
        RECT 71.850 153.980 72.150 154.980 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER Metal5 ;
        RECT 68.010 153.980 68.310 154.980 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER Metal5 ;
        RECT 64.170 153.980 64.470 154.980 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER Metal5 ;
        RECT 60.330 153.980 60.630 154.980 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER Metal5 ;
        RECT 117.930 153.980 118.230 154.980 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER Metal5 ;
        RECT 114.090 153.980 114.390 154.980 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER Metal5 ;
        RECT 110.250 153.980 110.550 154.980 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER Metal5 ;
        RECT 106.410 153.980 106.710 154.980 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER Metal5 ;
        RECT 102.570 153.980 102.870 154.980 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER Metal5 ;
        RECT 98.730 153.980 99.030 154.980 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER Metal5 ;
        RECT 94.890 153.980 95.190 154.980 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER Metal5 ;
        RECT 91.050 153.980 91.350 154.980 ;
    END
  END uo_out[7]
  PIN VGND
    PORT
      LAYER Metal5 ;
        RECT 16.000 0.000 18.200 152.980 ;
    END
  END VGND
  PIN VPWR
    PORT
      LAYER Metal5 ;
        RECT 20.000 0.000 22.200 152.980 ;
    END
  END VPWR
  OBS
      LAYER TopMetal2 ;
        RECT 0.000 153.730 11.060 154.980 ;
      LAYER TopMetal2 ;
        RECT 11.060 153.730 202.080 154.980 ;
      LAYER TopMetal2 ;
        RECT 0.000 149.260 3.295 153.730 ;
      LAYER TopMetal2 ;
        RECT 3.295 149.260 202.080 153.730 ;
      LAYER TopMetal2 ;
        RECT 0.000 148.000 11.060 149.260 ;
      LAYER TopMetal2 ;
        RECT 11.060 148.000 202.080 149.260 ;
      LAYER TopMetal2 ;
        RECT 0.000 146.000 202.080 148.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 129.000 202.080 146.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 127.000 202.080 129.000 ;
        RECT 0.000 126.205 11.060 127.000 ;
      LAYER TopMetal2 ;
        RECT 11.060 126.205 202.080 127.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 121.735 3.295 126.205 ;
      LAYER TopMetal2 ;
        RECT 3.295 121.735 202.080 126.205 ;
      LAYER TopMetal2 ;
        RECT 0.000 119.735 11.060 121.735 ;
      LAYER TopMetal2 ;
        RECT 11.060 119.735 202.080 121.735 ;
      LAYER TopMetal2 ;
        RECT 0.000 115.265 3.295 119.735 ;
      LAYER TopMetal2 ;
        RECT 3.295 115.265 202.080 119.735 ;
      LAYER TopMetal2 ;
        RECT 0.000 113.265 11.060 115.265 ;
      LAYER TopMetal2 ;
        RECT 11.060 113.265 202.080 115.265 ;
      LAYER TopMetal2 ;
        RECT 0.000 108.795 3.295 113.265 ;
      LAYER TopMetal2 ;
        RECT 3.295 108.795 202.080 113.265 ;
      LAYER TopMetal2 ;
        RECT 0.000 108.000 11.060 108.795 ;
      LAYER TopMetal2 ;
        RECT 11.060 108.000 202.080 108.795 ;
      LAYER TopMetal2 ;
        RECT 0.000 106.000 202.080 108.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 89.000 202.080 106.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 87.000 202.080 89.000 ;
        RECT 0.000 86.205 11.060 87.000 ;
      LAYER TopMetal2 ;
        RECT 11.060 86.205 202.080 87.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 81.735 3.295 86.205 ;
      LAYER TopMetal2 ;
        RECT 3.295 81.735 202.080 86.205 ;
      LAYER TopMetal2 ;
        RECT 0.000 79.735 11.060 81.735 ;
      LAYER TopMetal2 ;
        RECT 11.060 79.735 202.080 81.735 ;
      LAYER TopMetal2 ;
        RECT 0.000 75.265 3.295 79.735 ;
      LAYER TopMetal2 ;
        RECT 3.295 75.265 202.080 79.735 ;
      LAYER TopMetal2 ;
        RECT 0.000 73.265 11.060 75.265 ;
      LAYER TopMetal2 ;
        RECT 11.060 73.265 202.080 75.265 ;
      LAYER TopMetal2 ;
        RECT 0.000 68.795 3.295 73.265 ;
      LAYER TopMetal2 ;
        RECT 3.295 68.795 202.080 73.265 ;
      LAYER TopMetal2 ;
        RECT 0.000 68.000 11.060 68.795 ;
      LAYER TopMetal2 ;
        RECT 11.060 68.000 202.080 68.795 ;
      LAYER TopMetal2 ;
        RECT 0.000 66.000 202.080 68.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 49.000 202.080 66.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 47.000 202.080 49.000 ;
        RECT 0.000 46.205 11.060 47.000 ;
      LAYER TopMetal2 ;
        RECT 11.060 46.205 202.080 47.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 41.735 3.295 46.205 ;
      LAYER TopMetal2 ;
        RECT 3.295 41.735 202.080 46.205 ;
      LAYER TopMetal2 ;
        RECT 0.000 39.735 11.060 41.735 ;
      LAYER TopMetal2 ;
        RECT 11.060 39.735 202.080 41.735 ;
      LAYER TopMetal2 ;
        RECT 0.000 35.265 3.295 39.735 ;
      LAYER TopMetal2 ;
        RECT 3.295 35.265 202.080 39.735 ;
      LAYER TopMetal2 ;
        RECT 0.000 33.265 11.060 35.265 ;
      LAYER TopMetal2 ;
        RECT 11.060 33.265 202.080 35.265 ;
      LAYER TopMetal2 ;
        RECT 0.000 28.795 3.295 33.265 ;
      LAYER TopMetal2 ;
        RECT 3.295 28.795 202.080 33.265 ;
      LAYER TopMetal2 ;
        RECT 0.000 28.000 11.060 28.795 ;
      LAYER TopMetal2 ;
        RECT 11.060 28.000 202.080 28.795 ;
      LAYER TopMetal2 ;
        RECT 0.000 26.000 202.080 28.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 9.000 202.080 26.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 7.000 202.080 9.000 ;
        RECT 0.000 5.730 11.060 7.000 ;
      LAYER TopMetal2 ;
        RECT 11.060 5.730 202.080 7.000 ;
      LAYER TopMetal2 ;
        RECT 0.000 1.260 3.295 5.730 ;
      LAYER TopMetal2 ;
        RECT 3.295 1.260 202.080 5.730 ;
      LAYER TopMetal2 ;
        RECT 0.000 0.000 11.060 1.260 ;
      LAYER TopMetal2 ;
        RECT 11.060 0.000 202.080 1.260 ;
  END
END tt_um_htfab_yadge
END LIBRARY

